
//Global defines

`define AHB_ADDR_WIDTH 32
`define AHB_DATA_WIDTH 32
`define NONSEQ 2'b10
`define IDLE 2'b00
`define OKAY   	2'b00
`define ERROR   2'b01
