/*
 Licensed under the Apache License, Version 2.0 (the "License");         
 you may not use this file except in compliance with the License.        
 You may obtain a copy of the License at                                 
                                                                         
     http://www.apache.org/licenses/LICENSE-2.0                          
                                                                         
  Unless required by applicable law or agreed to in writing, software    
 distributed under the License is distributed on an "AS IS" BASIS,       
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and     
 limitations under the License.      
*/

//==============================================================||
// File Name: 		en_cnt.v				||
// Author:    		Kitty Wang				||
// Description: 						||
//	      		en count			       	|| 
// History:   							||
//                      2019/1/22 				||
//                      First version				||
//===============================================================


module en_cnt (
input wire clk,
input wire rstn,
input wire en,
output reg [31:0] cnt
);

always @ (posedge clk or negedge rstn)
begin
	if(!rstn)
	begin
		cnt <= 0;
	end
	else
	begin 
		if(en)
		begin
			cnt <= cnt + 1;
		end
	end
end

endmodule
