//`define RISCV
//`define ZEPHYR
`define ZEPHYR_PHIL
//`define ZEPHYR_SYNC
//`define INT_TEST
//`define PG_TEST

